library verilog;
use verilog.vl_types.all;
entity MuxComportamental_8_1_vlg_vec_tst is
end MuxComportamental_8_1_vlg_vec_tst;
