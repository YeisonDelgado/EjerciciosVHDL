library verilog;
use verilog.vl_types.all;
entity Decodificador_4_2_vlg_check_tst is
    port(
        f               : in     vl_logic_vector(1 downto 0);
        sampler_rx      : in     vl_logic
    );
end Decodificador_4_2_vlg_check_tst;
