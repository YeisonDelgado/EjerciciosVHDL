library verilog;
use verilog.vl_types.all;
entity Decodificador_4_2_vlg_vec_tst is
end Decodificador_4_2_vlg_vec_tst;
