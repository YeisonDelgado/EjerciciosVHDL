library verilog;
use verilog.vl_types.all;
entity Ejercicio2_vlg_vec_tst is
end Ejercicio2_vlg_vec_tst;
