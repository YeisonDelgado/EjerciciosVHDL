library verilog;
use verilog.vl_types.all;
entity MuxComportamental_8_1_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MuxComportamental_8_1_vlg_check_tst;
